module one_to_four_Dmux(
    input 
);
    
endmodule